module ALU(
input[3:0] A,
input[3:0] B,
input[2:0] OpCode,
output reg[7:0] Result,
output reg Zero,
output reg Carry
);

always @(*) begin
Zero = 0;
Carry = 0;
case(OpCode)
3'b000: Result = A + B;
3'b001: Result = A - B;
3'b010: Result = A*B;
3'b011: Result = B!=0 ? A/B : 8'b0;
default: Result = 8'b0;
endcase
if (Result == 8'b0)
Zero = 1'b1;
if ((OpCode == 3'b000)&&(((A==4'b1111)&&(B>4'b0000))||((B == 4'b1111)&&(A>4'b0000))))
Carry = 1'b1;
end
endmodule


